library verilog;
use verilog.vl_types.all;
entity ALSU_tb is
end ALSU_tb;
